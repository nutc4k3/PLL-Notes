.include sky130nm.lib
.include PFD.spice

XX1 Ref_Clk Up Down Clk2 GND VDD PFD

v1 VDD GND 1.8v

v2 Ref_Clk GND PULSE 0 1.8v 0 6p 6p 40n 80n

v3 Clk2 GND PULSE 0 1.8v 1n 6p 6p 40n 80n

.control 
tran 0.1n 5u
plot v(Up) v(Down)+2 v(Ref_Clk)+4 v(Clk2)+6
.endc

.end